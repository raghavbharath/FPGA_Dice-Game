library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_ARITH.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;
library lpm;
use lpm.lpm_components.all;

entity lab5_part4 is 
port (clk: in std_logic;
		button: in std_logic;
		display1: out std_logic_vector(0 to 6);
		display2: out std_logic_vector(0 to 6);
		display3: out std_logic_vector(0 to 6);
		display4: out std_logic_vector(0 to 6);
		die_value1: out std_logic_vector(2 downto 0);
		die_value2: out std_logic_vector(2 downto 0);
		die_value3: out std_logic_vector(2 downto 0);
		die_value4: out std_logic_vector(2 downto 0)
		);
		
end lab5_part4;

architecture structural of lab5_part4 is 

component lab5_part3 
port (pulse: in std_logic;
		die: out std_logic_vector(0 to 6);
		die_val: out std_logic_vector(2 downto 0));
		
end component;


signal clkb, clk1, clk2, clk3, clk4: std_logic;

begin 

	clkb <= clk and (not button);
	
	delay1: lpm_counter 
	generic map(lpm_width=>4) 
	port map (clock=>clkb, cout=> clk1);
	delay2: lpm_counter 
	generic map(lpm_width=>5) 
	port map (clock=>clkb, cout=> clk2);
	delay3: lpm_counter 
	generic map(lpm_width=>6) 
	port map (clock=>clkb, cout=> clk3);
	delay4: lpm_counter 
	generic map(lpm_width=>7) 
	port map (clock=>clkb, cout=> clk4);
	
	die1: lab5_part3 port map(die_val => die_value1,pulse => clk1, die(0 to 6) => display1(0 to 6));
	die2: lab5_part3 port map(die_val => die_value2,pulse => clk2, die(0 to 6) => display2(0 to 6));
	die3: lab5_part3 port map(die_val => die_value3,pulse => clk3, die(0 to 6) => display3(0 to 6));
	die4: lab5_part3 port map(die_val => die_value4,pulse => clk4, die(0 to 6) => display4(0 to 6));
	
end structural;

	